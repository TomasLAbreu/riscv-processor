
// ============================================================================
// riscv pipeline processor
// ============================================================================
//
// follows 5 cycle stages through a pipeline:
//    if    instruction fetch
//    id    instruction decode
//    ex    execute
//    mem   access data memory
//    wb    writeback
//
// ============================================================================

//------------------------------------------------------------------------------
module riscv
//------------------------------------------------------------------------------
#(
  parameter MP_DATA_WIDTH = 32,
  parameter MP_ADDR_WIDTH = 5,
  parameter MP_ENDIANESS = `RISCV_BIG_ENDIAN
)
(
	//TODO: parameterize instr* and PC
	//TODO: change rst to rstn
  input wire                        iclk,
  input wire                        irst,

  // Instruction memory
  input  wire [31:0]                iinstr, // Instruction
  output wire [31:0]                opc,    // Program counter

  // Data memory
  output wire [31:0]                odmem_addr,
  output wire [1:0]                 odmem_wr_be,
  output wire                       odmem_wr_en,
  output wire [MP_DATA_WIDTH-1 : 0] odmem_wr_data,
  input  wire [MP_DATA_WIDTH-1 : 0] idmem_rd_data
);
//------------------------------------------------------------------------------

  // ------ controler outputs
  wire [2:0] wctrl_rd_wr_data_src;
  wire wctrl_alu_src;

  wire wctrl_rd_wr_en_2d;
  wire wctrl_rd_wr_en_1d;

  wire wctrl_pc_result_src;
  wire [2:0] wctrl_imm_src;
  wire [3:0] wctrl_alu_ctrl;
  wire wctrl_result_srcb0;

  // ------ datapath outputs
  wire [4:0] wdp_rs1;
  wire [4:0] wdp_rs2;
  wire [4:0] wdp_rs1_1d;
  wire [4:0] wdp_rs2_1d;
  wire [4:0] wdp_rd;
  wire wctrl_pc_src;

  wire [4:0] wdp_rd_1d;
  wire [4:0] wdp_rd_2d;

  wire [31:0] wdp_instr;

  // ALU flags
  wire wdp_alu_zero;
  wire wdp_alu_ovfl;
  wire wdp_alu_carry;
  wire wdp_alu_neg;

  // ------ hazard unit flags
  wire [1:0] whazard_forward_alu_src_a;
  wire [1:0] whazard_forward_alu_src_b;
  wire whazard_stall_if;
  wire whazard_stall_id;
  wire whazard_flush_id;
  wire whazard_flush_ex;

  wire [6:0] wop;
  wire [2:0] wfunct3;
  wire wfunct7b5;

  assign wop = wdp_instr[6:0];
  assign wfunct3 = wdp_instr[14:12];
  assign wfunct7b5 = wdp_instr[30];

  riscv_ctrl u_ctrl (
    .iclk           (iclk),
    .irst           (irst),
    .iflush_e       (whazard_flush_ex),
    .iop            (wop),
    .ifunct3        (wfunct3),
    .ifunct7b5      (wfunct7b5),
    .oalu_src       (wctrl_alu_src),
    .oalu_ctrl      (wctrl_alu_ctrl),
    .ialu_zero      (wdp_alu_zero),
    .ialu_ovfl      (wdp_alu_ovfl),
    .ialu_carry     (wdp_alu_carry),
    .ialu_neg       (wdp_alu_neg),
    .oresult_src_2d (wctrl_rd_wr_data_src),
    .oresult_srcb0  (wctrl_result_srcb0),
    .odmem_wr_en    (odmem_wr_en),
    .ord_wr_en_1d   (wctrl_rd_wr_en_1d),
    .ord_wr_en_2d   (wctrl_rd_wr_en_2d),
    .opc_src        (wctrl_pc_src),
    .opc_result_src (wctrl_pc_result_src),
    .oimm_src       (wctrl_imm_src)
  );

  riscv_dp #(
    .MP_DATA_WIDTH (MP_DATA_WIDTH),
    .MP_ADDR_WIDTH (MP_ADDR_WIDTH),
    .MP_ENDIANESS  (MP_ENDIANESS)
  ) u_datapath (
    .iclk               (iclk),
    .irst               (irst),
    .iforward_alu_src_a (whazard_forward_alu_src_a),
    .iforward_alu_src_b (whazard_forward_alu_src_b),
    .istall_f           (whazard_stall_if),
    .istall_d           (whazard_stall_id),
    .iflush_d           (whazard_flush_id),
    .iflush_e           (whazard_flush_ex),
    .iinstr_nxt         (iinstr),
    .oinstr             (wdp_instr),
    .ipc_src            (wctrl_pc_src),
    .ipc_result_src     (wctrl_pc_result_src),
    .opc                (opc),
    .iimm_src           (wctrl_imm_src),
    .ors1               (wdp_rs1),
    .ors1_1d            (wdp_rs1_1d),
    .ors2               (wdp_rs2),
    .ors2_1d            (wdp_rs2_1d),
    .ird_wr_en          (wctrl_rd_wr_en_2d),
    .ird_wr_data_src    (wctrl_rd_wr_data_src), // TODO: rename this?
    .ord                (wdp_rd),
    .ord_1d             (wdp_rd_1d),
    .ord_2d             (wdp_rd_2d),
    .ialu_ctrl          (wctrl_alu_ctrl),
    .ialu_src           (wctrl_alu_src),
    .oalu_result        (odmem_addr),
    .oalu_zero          (wdp_alu_zero),
    .oalu_ovfl          (wdp_alu_ovfl),
    .oalu_carry         (wdp_alu_carry),
    .oalu_neg           (wdp_alu_neg),
    .odmem_wr_data      (odmem_wr_data),
    .idmem_rd_data      (idmem_rd_data),
    .odmem_wr_be        (odmem_wr_be)
  );

	riscv_hazard_unit u_hazard_unit (
    .ipc_src            (wctrl_pc_src),
    .iresult_srcb0      (wctrl_result_srcb0),
    .irs1               (wdp_rs1),
    .irs1_1d            (wdp_rs1_1d),
    .irs2               (wdp_rs2),
    .irs2_1d            (wdp_rs2_1d),
    .ird                (wdp_rd),
    .ird_1d             (wdp_rd_1d),
    .ird_2d             (wdp_rd_2d),
    .ird_wr_en_1d        (wctrl_rd_wr_en_1d),
    .ird_wr_en_2d         (wctrl_rd_wr_en_2d),
    .oforward_alu_src_a (whazard_forward_alu_src_a),
    .oforward_alu_src_b (whazard_forward_alu_src_b),
    .ostall_f          (whazard_stall_if),
    .ostall_d          (whazard_stall_id),
    .oflush_d          (whazard_flush_id),
    .oflush_e          (whazard_flush_ex)
	);

endmodule
